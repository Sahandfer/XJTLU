* C:\Users\sahand.sabour16\Desktop\Schematic2.sch

* Schematics Version 9.1 - Web Update 1
* Thu Nov 08 16:33:42 2018



** Analysis setup **
.DC LIN V_V3 -9 9 1 
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic2.net"
.INC "Schematic2.als"


.probe


.END
